****** Analysis Section ******
.TRAN 10p 10n

******************************