****** Analysis Section ******
.TRAN 100p 2.6u

******************************
