*DEFINICION DE PARAMETROS

.PARAM Vdd1=1.1
.PARAM Tech = 32e-9
.PARAM UNIT_W = '2*Tech'
.PARAM UNIT_L = Tech