****** Analysis Section ******
.TRAN 100p 1.2u

******************************
