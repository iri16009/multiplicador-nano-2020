****** Analysis Section ******
.TRAN 10p 48.5n

******************************